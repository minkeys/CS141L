module testbench();
// Declare inputs as regs and outputs as wires
reg [7:0] startAddress;
reg clk;
reg start;

// wire [7:0] currentpc;

// Initialize all variables
initial begin        
	clk = 1;       // initial value of clock
	start = 1;  	// initial value of reset
	startAddress = 0;     // initial value of wenable
	
	#10  start = 1;    // use reset to set pc to 0
	#10  start = 0;    // end of reset pulse.
	#10      // wait a cycle, make sure the PC doesn't change
	#10
	#10  
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10  start = 0;

 end

// Clock generator
always begin
   #1  clk = ~clk; // Toggle clock every 5 ticks
						// this makes the clock cycle 10 ticks
end

// the following creates an instance of our program_counter register.
//   I copied this code verbatim from the walkthough.v that was
//   generated by Quartus when I created the .v file from the .bdf.


busmux_0	b2v_bm1(
	.sel(SYNTHESIZED_WIRE_26),
	.dataa(SYNTHESIZED_WIRE_1),
	.datab(SYNTHESIZED_WIRE_2),
	.result(SYNTHESIZED_WIRE_16));


busmux_1	b2v_bm2(
	.sel(SYNTHESIZED_WIRE_3),
	.dataa(SYNTHESIZED_WIRE_4),
	.datab(SYNTHESIZED_WIRE_5),
	.result(SYNTHESIZED_WIRE_10));


instructionROM	b2v_inst(
	.program_counter(SYNTHESIZED_WIRE_27),
	.branchFlag(SYNTHESIZED_WIRE_22),
	.labelFlag(SYNTHESIZED_WIRE_26),
	.immediateFlag(SYNTHESIZED_WIRE_3),
	.signFlag(SYNTHESIZED_WIRE_8),
	.haltFlag(SYNTHESIZED_WIRE_7),
	.instruction(instruction),
	.labelValue(SYNTHESIZED_WIRE_1),
	.opcode(SYNTHESIZED_WIRE_11),
	.rd(SYNTHESIZED_WIRE_18),
	.rs(SYNTHESIZED_WIRE_19),
	.rt(SYNTHESIZED_WIRE_20),
	.value(SYNTHESIZED_WIRE_4));


\21mux 	b2v_inst27(
	.S(SYNTHESIZED_WIRE_7),
	
	.A(clk),
	.Y(SYNTHESIZED_WIRE_28));


alu	b2v_inst29(
	.signFlag(SYNTHESIZED_WIRE_8),
	.input0(SYNTHESIZED_WIRE_9),
	.input1(SYNTHESIZED_WIRE_10),
	.opcode(SYNTHESIZED_WIRE_11),
	.overflowFlag(SYNTHESIZED_WIRE_15),
	.lessThanFlag(SYNTHESIZED_WIRE_23),
	.overflow(SYNTHESIZED_WIRE_17),
	.result(SYNTHESIZED_WIRE_2));


regfile32x8	b2v_inst9(
	.clock(SYNTHESIZED_WIRE_28),
	.regwriteFlag(SYNTHESIZED_WIRE_26),
	.labelFlag(SYNTHESIZED_WIRE_26),
	.overflowFlag(SYNTHESIZED_WIRE_15),
	.dataIn(SYNTHESIZED_WIRE_16),
	.overflowIn(SYNTHESIZED_WIRE_17),
	.rd(SYNTHESIZED_WIRE_18),
	.rs(SYNTHESIZED_WIRE_19),
	.rt(SYNTHESIZED_WIRE_20),
	.branchAddress(SYNTHESIZED_WIRE_25),
	.regA(SYNTHESIZED_WIRE_9),
	.regB(SYNTHESIZED_WIRE_5));


program_counter_logic	b2v_pcl(
	.clk(SYNTHESIZED_WIRE_28),
	.start(start),
	.branch(SYNTHESIZED_WIRE_22),
	.taken(SYNTHESIZED_WIRE_23),
	.inputPC(SYNTHESIZED_WIRE_27),
	.startAddress(startAddress),
	.target(SYNTHESIZED_WIRE_25),
	.outputPC(SYNTHESIZED_WIRE_27));



endmodule