module testbenchdup();
// Declare inputs as regs and outputs as wires
reg [7:0] inp0;
reg [7:0] inp1;
reg [3:0] opc;
reg clk;
reg signfl;



// wire [7:0] currentpc;

// Initialize all variables
initial begin        
	clk = 1;       // initial value of clock

	
	#10      // wait a cycle, make sure the PC doesn't change
	#10	inp0 = 2; inp1 = 4; opc = 0; signfl = 1;
	#10
	#10	inp0 = 1; inp1 = 3; opc = 1; signfl = 1;
	#10
	#10	inp0 = 23; inp1 = 32; opc = 2; signfl = 1;
	#10
	#10	inp0 = 23; inp1 = -32; opc = 2; signfl = 1;
	#10
	#10	inp0 = 5; inp1 = 7; opc = 3; signfl = 1;
	#10
	#10	inp0 = 6; inp1 = 8; opc = 4; signfl = 1;
	#10   
	#10	inp0 = 23; inp1 = 32; opc = 2; signfl = 1;
	#10
	#10	inp0 = 23; inp1 = 32; opc = 2; signfl = 1;
	#10
	#10	inp0 = 23; inp1 = 32; opc = 2; signfl = 1;
	#10
	#10	inp0 = 23; inp1 = 32; opc = 2; signfl = 1;
	#10
	#10	inp0 = 23; inp1 = 32; opc = 2; signfl = 1;
	#10
	#10	inp0 = 23; inp1 = 32; opc = 2; signfl = 1;
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10
	#10 inp0 = 23; inp1 = 32; opc = 2; signfl = 1;

 end

// Clock generator
always begin
   #5  clk = ~clk; // Toggle clock every 5 ticks
						// this makes the clock cycle 10 ticks
end

// the following creates an instance of our program_counter register.
//   I copied this code verbatim from the walkthough.v that was
//   generated by Quartus when I created the .v file from the .bdf.


alu	b2v_inst(
	.signFlag(signfl),
	.input0(inp0),
	.input1(inp1),
	.opcode(opc),
	.overflowFlag(ovfl),
	.lessThanFlag(ltfl),
	.overflow(SYNTHESIZED_WIRE_7),
	.result(res));

endmodule